BZh91AY&SY���� )߀Ryg������?���`{�@� $  D
G2h�14�@��`�M4 a2dшbi���4�&&�h �dɣ��i�0LM4��j��4 ѐ  �  � "���O�F��Jz���3S=S�i��z���B@6�ړĞ&�&��M2z��>ԉ���A�R�	��pO�U�$�I /�
�� �$����ol�&yt�W�}<�<{�����ܰWHg*$�(9X�Q�@6�r�?~��|-! ��NJY
y���/�\��ur�B�_Vߚ���2�X�-�5G�����yM=!�M�ˌ��T������L�wʃP�yxp+X]���9���ۉ� _Y@���r�͆Ώ1��1�����܆�45w���>��y��U�Q�s+ �оC\����b�-kI|d	��>K<����+�!���N]۬S$j��X�Y��DlC�o()	1b���xvdB�鿱fy�Z"C�D�ļ�� x��`�х5�ۛe��.��X�l{��ޖpMd�I�t*���zw逶��j-ߙ�C�����_KM�f�}4�.����e�(����;N��<q�$>�
$�$�I$�IOBJ�)3�{֩߹|�6�}��8�$$�D��B�AA�X,����\1Z�!�@����/�K6[�4U����k��CS�C9Ls��(V7�%�JS�g�vY5Y�@�)b�Be-����	$��,�qu��|�~�[\��y����ԛ��-`����8��+�����b@�hs/o絥��~\�VD�5��;Ͽ������}�˦����
SC��Rd�l��>�٣%YA�y���P�'�X>K�>��X&!�d[�D���T1KD�2�bD��~'�O߇�9;l/Z<����ִloc���.���#�c�'����}�����c�9`'ݤ��=�F���Dvc���ޯ�\	��{K�E������/��imz}o���I��+��%�/)����ǌ��#��J�n,0 \�
~J���d�`�ek���
 n(�!A`,�l)5�m/�r��!$���p<I٪$ˈL�M���)N��Ʀ*pB���B�e�څ��@\�����B'��Rw�|�t����;P)MG0{p�$b��CR�;��H
�XRpR��.F���+1��}=~ 3��gws���ޠ����� h<��	����[�T��z��	 n]�9�+���f� qӚ��o]����Cԃ�f�;B5B���0�!�4_@㩑aSx(x}4�� [�%F�,|������y�~P灚�HE�� �/���
=� Tٰ�A
�ZSA�b�`F�r 2�j��H(
��W?��B���Ma�h�,P��yN��w�m��εL���H�C�� ��?Z߳�hq���9��$ [�η޻¥�!�
H@l�t��k�u�7����(lR�/�$*��j��6�;ĳ\[�0�A �BL"���F-���~���t{�d��\ܼ���ON̐ؼ2�CB�B��5�LvV���d#��ʡ��ۗ��`��0)`�~%.����\ٷ���9Α"2"d�P��sU�:s���N��q�@��gn}@�R��ɹ��W���<'7�$��B �{' HT�q��eN��-�%�]�\�GPu�٘g�ݡ���ٴ����8�> !b��rD^�j�P���"�(HI�ct 