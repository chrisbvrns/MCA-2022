BZh91AY&SY�v�� �߀Ryg������?���`�P �44 
	"M����  � 4 �h�L��M`&i�L� �2hb14`��@	��24	SS@�z��@4hѠi�h  �dɡ��рFa `&�4��$H  S  �$4�S�mCF���bD��4�)(B	� �$�SB��1�x�� $.��zZO��*"�Ln���M
Ig��c����@4�� D� V@��Hb�(J��?�fƕ���[��Ǫ��>5��K�ո$���/&R���20޾DL�ѽ� �J����~���fc���j"�m� �b���)g7�{)k�[;����a�_,���`�ĉ�
bJHsB ��Hڋ�H�w��F%���4�cWWN��K�^�����(�H�!.OɆƓsiC�&_���B��|-A&�lZsh�t�,���M�0x:�S�(�&H}fP���U!)]�I����"c�֡;4X\XA�b�а+5`R����l8`���`�����m���C�V�^Z\к�a%/�Ռ�Ln�r�pwApH$h�IL)��(��3�$\�d�Nf/$2�$)�S"�A�����'PakB�
8��Km����_|%��l�Z�Yff�K��8��#���`�̈́����w���/�TG�b�y�����vX��Ai 8���,�fE������k>=�vLЕE>r�Q��/XlFv^�zlg�h��"@��;сV&�`�	H=���v�<��xs)��h�%zI����h�������I_�nx���F7� �iD���l�>��Ȁ�"�G�)i �G��X�"'9϶s�l���J��^��kcV�o3�h�ē�C��3���Ia9��.ٕ�T2'M@"*,"�d��o�C w��>��,�&8�t]���������>�9
��~�=�N���(U/��
y'i�~L>f��1�j���PG`HcL}tޏ���F��$��%3�Li��%4�qb��z����n�P���A)`�:4��q
����&��zG k�XRpw�h]A�p���4r6���SC/
� u�R��h�i� �X��p.*HH�
���B?
�E�j���)LԁH���5w�*�b�PJj�}���APC��d5'
��$�n�H�Uw"��L !CH���;j�a�⸹��J�A�
έ�� |؛�tp&�z��h9f6/?>4?�pi��9g�p1g��5�D��8-Kd���Hr[o9�1�Jm-���nnJȲJ���k�0��#a&�K=�U�JCuS��r��^��Bf(f�F z���J��f��(A.iϬ�����$����¾�L��WL�0L),G"��k7A��� ebL�fXX�4˒�\��ը����a�V�%��*Ĵ�GN�D���FƁ�����`dH[Qq�@���a�3#4i5���9��P��G���%�2T����/��������`�5�����]��BB�ڛP