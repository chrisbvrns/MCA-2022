BZh91AY&SY�� �_�Ryg������?���`�z�    J��OS�  a �4� �&M�&�L�bi��!�L�1M00&�#��M A)�UF@Ѧ��1 � q�&�CL	��14�@H�@F@�4���К�P��(�G�)0G�38�\|��&���5M
����[0��(�cd��g�Ƈ)�9��R��T5�Ym��1�1��@4�� D� + J�A$1l�%V�#X3cJ��\�������俾?�|=it[�;�'}
̓��"!�T-g4M���j��Z�������*:��Z���c���P	Y�d���墖�%����d��1bݯ��ZZm�.zC�Ȕ���hIQi��H]�Ӱ��d\wf��j�ժW.S����|Y�R(D,YB�Ndf�xNb�ư������x
I��A��8`����%�3f#iRA�b�v%b�
ͬq��y;I�+!�VcRƊ���H(�y�T-/��v%QDa3��6�f�9YR܄�ʪ����3�3�����W`�0���%p3��FS	)��]ϺV�w��C$2!�b��/�i[����MD�L��)١c$\�A��0(�]����m!���X�����u����N�!�v	�/Dw�J�F$H�FQ�`xD���G�k�����KNϑ�6�e���ӝJ���
�KϣI��^�xl7����huK8�É���/0W��}�d����gY�k�bV�{��A��q�#�z.m�63��� _1���p��JA���=���A��-ׇJ�����i�,�,Ns���Dִ��O�;hx��7��dO�kg����F$ ���$�:c�����e���"s��'>|+jЕ۸����#pe9���������3��t�6�<�_@P��`
�N��h!B��,@IIu� ;�`G�%x1�\��:�eh��<y1.)H{�{@�k��N�z
�>��X�݇�
��H�ʐ�Ԋ��F�4��ƛ����ch�D�xhS<	�0�D��� ;9#�o' ,�p�5��h/�/�D��\��>��R�T��ҷ1��5�,)>���=7�&)����J7�`(e�� Σ��[��$gBì!K��⤄� TG`�#�P��MCP0g�0cR!�� ^on�c��T��k���u�A��`d5'
���5��*�]Ȥ��EP�"&|;*���x�.e0R�A�
ήU� |07 �<�M���	�ߠl>nE>Z�=����F��������Z$$g�ԶL z3�m��p�J���C_[p��Fd�z�I�2��^��v��Is#�%44Ҁ���_��GAiw7��Й�2b�����E�,h#���
o�	��d��|�9�0�}oC%4���K�L),G"�����l 4U&l4�0G<˒�]*v����a���ëU��pbY�:�4����#���lG9�G#���L����7�)�ٸ7�����I}0T���0_�>��s�����L�4�rE8P���