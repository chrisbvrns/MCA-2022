BZh91AY&SY��  w_�Pyc���ߺ?���P��wq�$6��l����F�� �	��O	��!���h� ɣCL��4�"B512��)�i��4� � h2d�L&F@��M#4i�RM	�S�4�jOOe���i� ���)�����L<��̧x��J���3��q�5�GBh��mcJ�Ј ����XR��9���"l�<2��]cv���[h�b}rn��|�HU$e�a�S!��r�T���D$����3[5����x��l�%�	�C��K!	����Lɥˮ63������-&#Q�ЮШF%��f4)��-�ȶ1����m���d'b2l$U+2D��Y2�M��XJ��ժ*ɰrk{_�+�<��P���CF��*�iP f
�q��j�7��i�Qt�<����H�*��N1ș�V�Ǯ�<%��o0�H��;�4�(-	���'q�������zZ�zB���1$�[C�	9��}i�փ��������~(짝��$�q��Rc2�δ�I+6s3&����5U:�,��nS&������6�ݚ��u�LM�X�)K��(T��3�Qk
N$^l)۳C��+�K����Q �2${{�g�!F?M��u� F���-�7�>���h��G=L�Be�M'=c��p-
��iK#�b�������Ꮺ��7�T��;�n0�<N�H�J�S��v@d+�E��i��f$��A��$;�%�2F/ϐpI"����M@��H�-f��$�!e�i�!:%`�3��0�B��^��#��ޖ�k>���MN��P����{�!� q4��nm�b'!w�1!���1�8�M(��f��)�ٛ�b1��Ы׎8�h�l�9<k!+����D\-ҕH6�m8��a5���0&%��K��f&d�ۺ�����29�5���mP��MIMpN߄`A.�l.��]��BB�p 